interface dff_interface;
    logic clk;        // Clock signal
    logic rst;        // Reset signal
    logic din;        // Data input signal
    logic dout;       // Data output signal
endinterface : dff_interface
