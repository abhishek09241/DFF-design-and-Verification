package sim_dff_pkg;
			`include "transaction.sv"
			`include "generator.sv"
			`include "driver.sv"
			`include "monitor.sv"
			`include "scoreboard.sv"
			`include "environment.sv"
endpackage : sim_dff_pkg		