class scoreboard;
	transaction tr;					// Define a tansaction object
	transaction trref;				// Define a reference transaction object for comparison
	mailbox #(transaction) mbx;		// Create a mailbox to receive data from the driver
	mailbox	#(transaction) mbxref; 	// Create a mailbox to receive reference data from the generator
	event sconext;					// Event to signal completion of scoreboard work


	function new(mailbox #(transaction) mbx, mailbox #(transaction) mbxref);
		 	this.mbx 	= mbx;		// Initialize the mailbox for receiving data from the driver
		 	this.mbxref	= mbxref;	// Initialize the mailbox for receiving reference data from the generator		
	endfunction
	

	task run();
			forever
				begin
					mbx.get(tr);		// Get a transaction from the driver
					mbxref.get(trref);	// Get a reference transaction from the generator
					tr.display("SCO");	// Display the refenrece transaction information
					trref.display("REG");	// Display the reference transaction information
					if (tr.dout==trref.din)
						 begin
							$display("[SCO] : DATA MATCHED");		// Compare data and display the result
						end	
					else	
							$display("[SCO] : DATA MISMATCHED");
						$display("----------------------");
						->sconext; 		// Signal completion of scoreboard work
				end
	endtask : run	
endclass : scoreboard